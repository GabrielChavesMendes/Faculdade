module shift_register (
    input wire clk,
    input wire rst,
    input wire LD,
    input wire D,
    output reg [5:0] Q
);

always @(posedge clk or posedge rst) begin
    if (rst)
        Q <= 6'b0;
    else if (LD)
        Q[5:0] <= {D, Q[5:1]};
    else
        Q[5:0] <= {1'b0, Q[5:1]};
end

endmodule
